`ifndef AY_APB_DEF
`define AY_APB_DEF
    `ifndef AY_APB_MAX_DATA_WIDTH
        `define AY_APB_MAX_DATA_WIDTH 32
    `endif
    `ifndef AY_APB_MAX_ADDR_WIDTH
        `define AY_APB_MAX_ADDR_WIDTH 16
    `endif
`endif